module prf
import cpu_params::*;
(
    input   logic               clk,
    input   logic               rst,

    cdb_itf.prf                 cdb
);



endmodule
