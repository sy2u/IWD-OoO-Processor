module int_rs
import cpu_params::*;
(
    input   logic               clk,
    input   logic               rst,

    id_int_rs_itf.int_rs        from_id
);



endmodule
