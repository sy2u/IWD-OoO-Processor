module rat
import cpu_params::*;
(
    input   logic               clk,
    input   logic               rst,

    id_rat_itf.rat              from_id,
    cdb_itf.rat                 cdb
);



endmodule
