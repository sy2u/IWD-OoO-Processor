module free_list
import cpu_params::*;
(
    input   logic               clk,
    input   logic               rst,

    id_fl_itf.fl                from_id,
    rrf_fl_itf.fl               from_rrf
);



endmodule
