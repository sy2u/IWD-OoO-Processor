module fu_alu
import cpu_params::*;
(
    input   logic               clk,
    input   logic               rst,

    cdb_itf.fu                  cdb
);



endmodule
