module rrf
import cpu_params::*;
(
    input   logic               clk,
    input   logic               rst,

    rob_rrf_itf.rrf             from_rob,
    rrf_fl_itf.rrf              to_fl
);


endmodule
